$(header)

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
LIBRARY work;
USE work.types_pkg.ALL;

PACKAGE $(particle)_setup IS
$(eta_4)
$(phi_4)
$(eta_2_s)
$(phi_2_s)
$(eta_2_wsc)
$(phi_2_wsc)
-- $(control_2_wsc)
$(delta_eta)
$(delta_phi)
$(eta_1_s)
$(phi_1_s)
END $(particle)_setup;
-- dummy change --
-- dummy change --
-- dummy change --
